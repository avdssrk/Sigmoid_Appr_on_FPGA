`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   11:52:19 06/08/2023
// Design Name:   sigmoid1
// Module Name:   C:/Users/Pulak Mondal/Desktop/Shiva/Sigmoid_appr1/test_sigmoid.v
// Project Name:  Sigmoid_appr1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: sigmoid1
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test_sigmoid;

	// Inputs
	reg [15:0] in;

	// Outputs
	wire [15:0] out;

	// Instantiate the Unit Under Test (UUT)
	sigmoid1 uut (
		.in(in), 
		.out(out)
	);

	initial begin
		// Initialize Inputs
		in = 0;

		// Wait 100 ns for global reset to finish
		#100;
		
		in = 16'b1_1100_0000_0000_000;   //-4
		#100;
		
		in = 16'b1_1100_1000_0000_000;   //-3.5
		#100;
		
		in = 16'b1_1101_0000_0000_000;   //-3
		#100;
		
		in = 16'b1_1101_1000_0000_000;   //-2.5
		#100;
		
        in = 16'b1_1110_0000_0000_000;   //-2
		#100;
		
		in = 16'b1_1110_1000_0000_000;   //-1.5
		#100;
		
		in = 16'b1_1111_0000_0000_000;   //-1
		#100;
		
		in = 16'b1_1111_1000_0000_000;   //-0.5
		#100;
		
		in = 16'b00000_0000_0000_000;   //0
		#100;
		
		in = 16'b0_0000_1000_0000_000;   //0.5
		#100;
		
        in = 16'b0_0001_0000_0000_000;   //1
		#100;
        
		in = 16'b0_0001_1000_0000_000;   //1.5
		#100;
		
        in = 16'b0_0010_0000_0000_000;   //2
		#100;
        
		in = 16'b0_0010_1000_0000_000;   //2.5
		#100;
		
        in = 16'b0_0011_0000_0000_000;   //3
		#100;
		
		in = 16'b0_0011_1000_0000_000;   //3.5
		#100;
		
		in = 16'b0_0100_0000_0000_000;   //4
		#100;
		
		in = 16'b1_1111_0000_0000_000; //-1
		#100;
		
		in = 16'b1_1111_0001_1001_110; //-0.9
		#100;
		
		in = 16'b1_1111_0011_0011_010; //-0.8
		#100;
		
		in = 16'b1_1111_0100_1100_111; //-0.7
		#100;
		
		in = 16'b1_1111_0110_0110_100; //-0.6
		#100;
		
		in = 16'b1_1111_1000_0000_000; //-0.5
		#100;
		
		in = 16'b1_1111_1001_1001_101; //-0.4
		#100;
		
		in = 16'b1_1111_1011_0011_010; //-0.3
		#100;
		
		in = 16'b1_1111_1100_1100_111; //-0.2
		#100;
		
		in = 16'b1_1111_1110_0110_100; //-0.1
		#100;
		
		in = 16'b0_0000_0000_0000_000; //0
		#100;
		
		in = 16'b0_0000_0001_1001_100; //0.1
		#100;
		
		in = 16'b0_0000_0011_0100_000; //0.2
		#100;
		
		in = 16'b0_0000_0100_1100_110; //0.3 
		#100;
		
		in = 16'b0_0000_0110_0110_011; //0.4
		#100;
		
		in = 16'b0_0000_1000_0000_000; //0.5
		#100;
		
		in = 16'b0_0000_1001_1001_100; //0.6
		#100;
		
		in = 16'b0_0000_1011_0011_001; //0.7
		#100;
		
		in = 16'b0_0000_1100_1100_110; //0.8
		#100;
		
		in = 16'b0_0000_1110_0110_010; //0.9
		#100;
		
		in = 16'b0_0001_0000_0000_000; //1
		#100;
		
		
		// Add stimulus here

	end
      
endmodule

